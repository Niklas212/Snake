module main
/*
fn main() {
	mut snake:= Snake{}
	snake.field.set_food_random(snake)
	println(snake.get_map())
	snake.print()
}

fn (sn &Snake) print () {
	mut ret:=""
	m:=sn.get_map()
	for y in 0..sn.field.height {
		for x in 0..sn.field.width {
			ret+= match m[y][x] {
				1 {"@"}
				2 {"#"}
				3 {"*"}
				else {"."}
			}
		}
		ret+="\n"
	}
	
	println(ret)
}
*/